--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   02:21:54 04/08/2013
-- Design Name:   
-- Module Name:   /home/nilesh/Academics/cs288/Ping Pong/Paddle/debounce_Test.vhd
-- Project Name:  Paddle
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: debounce
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY debounce_Test IS
END debounce_Test;
 
ARCHITECTURE behavior OF debounce_Test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT debounce
    PORT(
         button : IN  std_logic;
         clk : IN  std_logic;
         outputLocked : OUT  std_logic;
         result : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal button : std_logic := '0';
   signal clk : std_logic := '0';

 	--Outputs
   signal outputLocked : std_logic;
   signal result : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: debounce PORT MAP (
          button => button,
          clk => clk,
          outputLocked => outputLocked,
          result => result
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		button<='1';
		wait for 1000 ns;
		button<='0';
		wait for 1000 ns;
		button<='1';
		
		
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
